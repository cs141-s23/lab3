module clk_divider
    (
        input logic clk_in, rst,
        output logic clk_out
    );

    // TODO: output one positive edge for every 100 million input positive edges

endmodule
