// define states
`define IDLE 4'b0000
`define SAMPLE_STATE1 4'b0001
`define SAMPLE_STATE2 4'b0010

// useful macros
`define LIGHT_RED 3'b001
`define LIGHT_YELLOW 3'b010
`define LIGHT_GREEN 3'b100

`define PED_NS 2'b10
`define PED_EW 2'b01
`define PED_BOTH 2'b11
`define PED_NEITHER 2'b00
