`include "tlc.svh"

module tlc_tb;

    // TODO: Your testbench here!

endmodule
